module Main #( parameter N = 32 )( input logic [N-1:0] x, output logic is_prime );
  assign is_prime = 1'b0;
endmodule